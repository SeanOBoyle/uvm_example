`ifndef DUT_SEQUENCE_LIST__SV
`define DUT_SEQUENCE_LIST__SV

// Base DUT Virtual Sequence
`include "dut_base_vseq.sv"

// Simple Test Sequence -- example
`include "dut_simple_vseq.sv"



`endif // DUT_SEQUENCE_LIST__SV