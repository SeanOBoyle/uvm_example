`ifndef HOST_SEQUENCE_LIST__SV
`define HOST_SEQUENCE_LIST__SV

`include "host_nominal_seq.sv"



`endif // HOST_SEQUENCE_LIST__SV