`ifndef  DUT_TEST_LIST__SV
 `define DUT_TEST_LIST__SV

// UVM/RUVM Packages
import uvm_pkg::*;

// Agents
import host_pkg::*;

`include "dut_test_base.sv"


`endif // DUT_TEST_LIST__SV
