`ifndef DUT_PKG__SV
`define DUT_PKG__SV

`include "uvm_macros.svh"
import uvm_pkg::*;

import host_pkg::*;


`include "dut_cfg.sv"
`include "dut_virtual_sequencer.sv"
`include "dut_env.sv"
`include "dut_sequence_list.sv"


`endif // DUT_PKG__SV